VGA_PLL_inst: VGA_PLL
port map(
          REFERENCECLK => ,
          PLLOUTCORE => ,
          PLLOUTGLOBAL => ,
          RESET => 
        );
