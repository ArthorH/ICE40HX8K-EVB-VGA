VGA_Clock_inst: VGA_Clock
port map(
          PACKAGEPIN => ,
          PLLOUTCORE => ,
          PLLOUTGLOBAL => ,
          RESET => 
        );
